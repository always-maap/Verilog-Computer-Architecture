module ALU(Control, A, B, Out, Zero);
    input [3:0] Control;
    input [31:0] A, B;
    
    output reg [31:0] Out;
    output Zero;
    
endmodule

module ALU_test;
    
endmodule